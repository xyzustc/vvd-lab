`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/04/01 07:18:46
// Design Name: 
// Module Name: alu
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module alu#(
    parameter WIDTH = 32
) (
    input [WIDTH-1:0] a,b,
    input [2:0] f,
    output [WIDTH-1:0] y,
    output z
);
reg [WIDTH-1:0] y_reg;
reg z_reg;

parameter f_plus = 3'b000;
parameter f_minus = 3'b001;
parameter f_and = 3'b010;
parameter f_or = 3'b011;
parameter f_xor = 3'b100;

assign y = y_reg;
assign z = z_reg;

always@(*) 
begin
    case(f)
        f_plus:     {y_reg,z_reg} = {a+b,0};
        f_minus:    {y_reg,z_reg} = {a-b,0};
        f_and:      {y_reg,z_reg} = {a&b,0};
        f_or:       {y_reg,z_reg} = {a|b,0};
        f_xor:      {y_reg,z_reg} = {a^b,0};
        default:    {y_reg,z_reg} = {0,1};
    endcase
end

//always@(*) 
//begin
////    if(f<=3'b100)   z_reg = 0;
////    else            z_reg = 1;
//    case(f)
//        f_plus:     z_reg = 0;
//        f_minus:    z_reg = 0;
//        f_and:      z_reg = 0;
//        f_or:       z_reg = 0;
//        f_xor:      z_reg = 0;
//        default:    z_reg = 1;
//    endcase
//end

endmodule

